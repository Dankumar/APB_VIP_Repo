
`include "uvm_macros.svh"
package apb_package;

 import uvm_pkg::*;
  `include "apb_define.sv"
  `include "apb_types.sv"
  `include "apb_env_cfg.sv"
  `include "apb_base_pkt.sv"
  `include "apb_sequencer.sv"
  `include "apb_sequence.sv"
  `include "apb_slave_monitor.sv"
  `include "apb_slave_driver.sv"
  `include "apb_master_monitor.sv"
  `include "apb_driver.sv"
  `include "apb_agent.sv"
  `include "apb_scoreboard.sv"
  `include "apb_env.sv"
endpackage
